decoder.sv

decode OPCODE {

    
}